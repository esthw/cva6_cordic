module sin_cos
    import ariane_pkg::*;
#(
    parameter config_pkg::cva6_cfg_t CVA6Cfg = config_pkg::cva6_cfg_empty
) (
    input  logic                             clk_i,
    input  logic                             rst_ni,
    input  logic                             flush_i,
    input  logic         [TRANS_ID_BITS-1:0] trans_id_i,
    input  logic                             valid_i,
    input  fu_op                             operation_i,
    input logic                       [63:0] fix64_in,
    output logic                      [63:0] fix64_out,
    output logic                             valid_o,
    output logic                             ready_o,
    output logic         [TRANS_ID_BITS-1:0] trans_id_o
);


    logic              [16:0] cnt;
    logic                     triangle_flag;
    logic signed       [63:0] sin;
    logic signed       [63:0] cos;
    logic signed       [63:0] data;
    fu_op                     operation, op0, op1, op2, op3, op4, op5, op6, op7, op8, op9, op10, op11, op12, op13, op14, op15, op16;


    logic signed 	    [63:0] x0=0,y0=0,z0=0;
    logic signed 	   	[63:0] x1=0,y1=0,z1=0;
    logic signed 	   	[63:0] x2=0,y2=0,z2=0;
    logic signed 	   	[63:0] x3=0,y3=0,z3=0;
    logic signed 	   	[63:0] x4=0,y4=0,z4=0;
    logic signed 	   	[63:0] x5=0,y5=0,z5=0;
    logic signed 	   	[63:0] x6=0,y6=0,z6=0;
    logic signed 	   	[63:0] x7=0,y7=0,z7=0;
    logic signed 	   	[63:0] x8=0,y8=0,z8=0;
    logic signed	   	[63:0] x9=0,y9=0,z9=0;
    logic signed 	   	[63:0] x10=0,y10=0,z10=0;
    logic signed 	   	[63:0] x11=0,y11=0,z11=0;
    logic signed 	   	[63:0] x12=0,y12=0,z12=0;
    logic signed 	   	[63:0] x13=0,y13=0,z13=0;
    logic signed 	   	[63:0] x14=0,y14=0,z14=0;
    logic signed 	   	[63:0] x15=0,y15=0,z15=0;
    logic signed 	   	[63:0] x16=0,y16=0,z16=0;

    logic signed        [63:0] result, result_q, result_d;
    logic               [TRANS_ID_BITS-1:0] id, id0, id1, id2, id3, id4, id5, id6, id7, id8, id9, id10, id11, id12, id13, id14, id15, id16;

// always_comb begin
//     if(valid_i)begin
//         data = fix64_in;
//     end
//     else begin
//         data = 'b0;
//     end

// end
assign data = valid_i ? fix64_in : 'b0 ;
assign operation = valid_i ? operation_i : 'b0 ;
assign id = valid_i ? trans_id_i : 'b0 ;
    

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x0    <= 64'b0; 						
		y0    <= 64'b0;
		z0    <= 64'b0;
        op0   <= 'b0;
        id0   <= 'b0;
	end
	else 
	begin
		x0    <= `k;
		y0    <=  64'd0;
		z0    <= data;
        op0   <= operation;
        id0   <= id;
	end

end


always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x1 <= 64'b0; 						
		y1 <= 64'b0;
		z1 <= 64'b0;
        op1   <= 'b0;
        id1 <= 'b0;
	end
	else
	begin
        op1   <= op0;
        id1   <= id0;
        if(z0[`sign_bit])
        begin
          x1 <= x0 + y0;
          y1 <= y0 - x0;
          z1 <= z0 + `rot0;
        end
        else
        begin
          x1 <= x0 - y0;
          y1 <= y0 + x0;
          z1 <= z0 - `rot0;
        end
	end

end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x2 <= 64'b0; 						
		y2 <= 64'b0;
		z2 <= 64'b0;
        op2<= 'b0;
        id2<= 'b0;
	end
	else 
	begin
        op2   <=  op1;
        id2   <=  id1;
	   if(z1[`sign_bit])
        begin
            x2 <= x1 + (y1 >>> 1);
            y2 <= y1 - (x1 >>> 1);
            z2 <= z1 + `rot1;
        end
        else
        begin
           x2 <= x1 - (y1 >>> 1);
           y2 <= y1 + (x1 >>> 1);
           z2 <= z1 - `rot1;
        end
    end
    
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x3 <= 64'b0; 						
		y3 <= 64'b0;
		z3 <= 64'b0;
        op3 <= 'b0;
	end
	else 
	begin
        op3   <= op2;
        id3 <= id2;
        if(z2[`sign_bit])
        begin
            x3 <= x2 + (y2 >>> 2);
            y3 <= y2 - (x2 >>> 2);
            z3 <= z2 + `rot2;
        end
        else
        begin
           x3 <= x2 - (y2 >>> 2);
           y3 <= y2 + (x2 >>> 2);
           z3 <= z2 - `rot2;
        end
    end
   
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x4 <= 64'b0; 						
		y4 <= 64'b0;
		z4 <= 64'b0;
        op4 <= 'b0;
	end
    else 
    begin
        op4   <= op3;
        id4 <= id3;
        if(z3[`sign_bit])
        begin
            x4 <= x3 + (y3 >>> 3);
            y4 <= y3 - (x3 >>> 3);
            z4 <= z3 + `rot3;
        end
        else
        begin
           x4 <= x3 - (y3 >>> 3);
           y4 <= y3 + (x3 >>> 3);
           z4 <= z3 - `rot3;
        end
    end
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x5 <= 64'b0; 						
		y5 <= 64'b0;
		z5 <= 64'b0;
        op5 <= 'b0 ;
        id5 <= 'b0 ;
	end
    else
    begin
        op5 <= op4;
        id5 <= id4;
        if(z4[`sign_bit])
        begin
            x5 <= x4 + (y4 >>> 4);
            y5 <= y4 - (x4 >>> 4);
            z5 <= z4 + `rot4;
        end
        else
        begin
           x5 <= x4 - (y4 >>> 4);
           y5 <= y4 + (x4 >>> 4);
           z5 <= z4 - `rot4;
        end
    end
    
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x6 <= 64'b0; 						
		y6 <= 64'b0;
		z6 <= 64'b0;
        op6 <= 'b0;
        id6 <= 'b0;
	end
    else
    begin
        op6 <= op5;
        id6 <= id5;
        if(z5[`sign_bit])
        begin
            x6 <= x5 + (y5 >>> 5);
            y6 <= y5 - (x5 >>> 5);
            z6 <= z5 + `rot5;
        end
        else
        begin
           x6 <= x5 - (y5 >>> 5);
           y6 <= y5 + (x5 >>> 5);
           z6 <= z5 - `rot5;
        end
    end
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x7 <= 64'b0; 						
		y7 <= 64'b0;
		z7 <= 64'b0;
        op7 <= 0 ;
        id7 <= 0 ;
	end
    else 
    begin
        op7 <= op6 ;
        id7 <= id6;
        if(z6[`sign_bit])
        begin
            x7 <= x6 + (y6 >>> 6);
            y7 <= y6 - (x6 >>> 6);
            z7 <= z6 + `rot6;
        end
        else
        begin
           x7 <= x6 - (y6 >>> 6);
           y7 <= y6 + (x6 >>> 6);
           z7 <= z6 - `rot6;
        end
    end
    
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x8 <= 64'b0; 						
		y8 <= 64'b0;
		z8 <= 64'b0;
        op8 <= 'b0 ;
        id8 <= 0;
	end
    else 
    begin
        op8 <= op7;
        id8 <= id7;
        if(z7[`sign_bit])
        begin
            x8 <= x7 + (y7 >>> 7);
            y8 <= y7 - (x7 >>> 7);
            z8 <= z7 + `rot7;
        end
        else
        begin
           x8 <= x7 - (y7 >>> 7);
           y8 <= y7 + (x7 >>> 7);
           z8 <= z7 - `rot7;
        end
    end
   
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x9 <= 64'b0; 						
		y9 <= 64'b0;
		z9 <= 64'b0;
        op9 <= 'b0;
        id9 <= 0;
	end
    else 
    begin
        op9 <= op8;
        id9 <= id8;
        if(z8[`sign_bit])
        begin
            x9 <= x8 + (y8 >>> 8);
            y9 <= y8 - (x8 >>> 8);
            z9 <= z8 + `rot8;
        end
        else
        begin
           x9 <= x8 - (y8 >>> 8);
           y9 <= y8 + (x8 >>> 8);
           z9 <= z8 - `rot8;
        end
    end
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x10 <= 64'b0; 						
		y10 <= 64'b0;
		z10 <= 64'b0;
        op10 <= 'b0 ;
        id10 <= 0;
	end
    else
    begin
        op10 <= op9 ;
        id10 <= id9 ;
        if(z9[`sign_bit])
        begin
            x10 <= x9 + (y9 >>> 9);
            y10 <= y9 - (x9 >>> 9);
            z10 <= z9 + `rot9;
        end
        else
        begin
           x10 <= x9 - (y9 >>> 9);
           y10 <= y9 + (x9 >>> 9);
           z10 <= z9 - `rot9;
        end
    end
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x11 <= 64'b0; 						
		y11 <= 64'b0;
		z11 <= 64'b0;
        op11 <= 'b0 ;
        id11 <= 0;
	end
    else 
    begin
        op11 <= op10;
        id11 <= id10;
        if(z10[`sign_bit])
        begin
            x11 <= x10 + (y10 >>> 10);
            y11 <= y10 - (x10 >>> 10);
            z11 <= z10 + `rot10;
        end
        else
        begin
           x11 <= x10 - (y10 >>> 10);
           y11 <= y10 + (x10 >>> 10);
           z11 <= z10 - `rot10;
        end
    end
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x12 <= 64'b0; 						
		y12 <= 64'b0;
		z12 <= 64'b0;
        op12 <= 'b0;
        id12 <= 0;
	end
    else 
    begin
        op12 <= op11 ;
        id12 <= id11 ;
        if(z11[`sign_bit])
        begin
            x12 <= x11 + (y11 >>> 11);
            y12 <= y11 - (x11 >>> 11);
            z12 <= z11 + `rot11;
        end
        else
        begin
           x12 <= x11 - (y11 >>> 11);
           y12 <= y11 + (x11 >>> 11);
           z12 <= z11 - `rot11;
        end
    end
    
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x13 <= 64'b0; 						
		y13 <= 64'b0;
		z13 <= 64'b0;
        op13 <= 'b0;
        id13 <= 0;
	end
    else
    begin
        op13 <= op12;
        id13 <= id12;
        if(z12[`sign_bit])
        begin
            x13 <= x12 + (y12 >>> 12);
            y13 <= y12 - (x12 >>> 12);
            z13 <= z12 + `rot12;
        end
        else
        begin
           x13 <= x12 - (y12 >>> 12);
           y13 <= y12 + (x12 >>> 12);
           z13 <= z12 - `rot12;
        end
    end
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x14 <= 64'b0; 						
		y14 <= 64'b0;
		z14 <= 64'b0;
        op14 <= 'b0;
        id14 <= 0;
	end
	else 
    begin
        op14 <= op13 ;
        id14 <= id13;
        if(z13[`sign_bit])
        begin
            x14 <= x13 + (y13 >>> 13);
            y14 <= y13 - (x13 >>> 13);
            z14 <= z13 + `rot13;
        end
        else
        begin
           x14 <= x13 - (y13 >>> 13);
           y14 <= y13 + (x13 >>> 13);
           z14 <= z13 - `rot13;
        end
    end
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x15 <= 64'b0; 						
		y15 <= 64'b0;
		z15 <= 64'b0;
        op15 <= 'b0 ;
        id15 <= 0;
	end
	else
    begin
        op15 <= op14;
        id15 <= id14;
        if(z14[`sign_bit])
        begin
            x15 <= x14 + (y14 >>> 14);
            y15 <= y14 - (x14 >>> 14);
            z15 <= z14 + `rot14;
        end
        else
        begin
           x15 <= x14 - (y14 >>> 14);
           y15 <= y14 + (x14 >>> 14);
           z15 <= z14 - `rot14;
        end
    end
end

always_ff @(posedge clk_i or negedge rst_ni)
begin
	if(!rst_ni || flush_i)
	begin
		x16 <= 64'b0; 						
		y16 <= 64'b0;
		z16 <= 64'b0;
        op16 <= 'b0 ;
        id16 <= 0;
		// cnt <= 0;
		// triangle_flag <= 1'b0;
		
	end
	else 
    begin
        op16 <= op15 ;
        id16 <= id15 ;
        if(z15[`sign_bit])
        begin
            x16 <= x15 + (y15 >>> 15);
            y16 <= y15 - (x15 >>> 15);
            z16 <= z15 + `rot15;
        end
        else
        begin
           x16 <= x15 - (y15 >>> 15);
           y16 <= y15 + (x15 >>> 15);
           z16 <= z15 - `rot15;
        end  
        
        // cnt <= cnt + 1;
        // if (cnt == 16)
        // begin
        //     triangle_flag <= 1'b1;
        //     trans_id_o <= trans_id_i; // ?
        // end
        // else
        // begin
        //     triangle_flag <= 1'b0;
        // end
            
    end
end


assign triangle_flag = (cnt[16]==1'b1) ? 1'b1 : 1'b0 ;
assign ready_o = 1'b1 ;  //?
// assign valid_o = ~flush_i && (operation_i inside {SIN, COS}) && triangle_flag ;
assign valid_o = ~flush_i && triangle_flag ;

// assign fix64_out = result_q;
// assign result = (op16==SIN) ? y16 : ((op16==COS) ? x16 : 'd0) ;
// assign result_d = valid_o ? result : result_q;
assign fix64_out = (op16==SIN) ? y16 : ((op16==COS) ? x16 : 'd0) ;

assign trans_id_o = id16 ;

//assign trans_id_o = trans_id_q;
//assign trans_id_d = valid_o ? trans_id_i : trans_id_q ;

always_ff @(posedge clk_i or negedge rst_ni)
begin
    if(!rst_ni || flush_i)
	begin
		cnt <= 0;
		// triangle_flag <= 1'b0;
        //result_q <= 0;
        //trans_id_q <= 0;
	end
    else begin
        // cnt[0] <= valid_i;
        // cnt <= {cnt[14:0], cnt[15]};
        cnt <= {cnt[15:0], valid_i};
        //result_q <= result_d;
        //trans_id_q <= trans_id_d;
    end
end


// always_comb begin

//     cos = x16; 						
// 	sin = y16;
   
    
//     if(operation_i == SIN)
//     begin
//         fix64_out = sin;  
//     end
//     else
//     begin
//          fix64_out = cos; 
//     end
// end
    
endmodule
